mudule a();



endmodule
