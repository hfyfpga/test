mudule a1();
input a;
input rst;

output ccpo;

endmodule
